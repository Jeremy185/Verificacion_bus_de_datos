`timescale 1ns / 1ps

module Ambiente(

    );
endmodule
